../xdc/psd_fpga_top.vh