../gpio/gpio_assigns.vh