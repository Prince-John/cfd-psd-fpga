`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07/25/2024 04:32:00 PM
// Design Name: 
// Module Name: psd_fpga_top
// Project Name: psd_fpga
// Target Devices: 
// Tool Versions: 
// Description: FPGA for PSD system
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

// %%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
// Include the top level module declaration
// DO NOT modify
// It is auto generated by the pin2xdc.tcl constraint generator
// %%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%

module psd_fpga_top(

`include    "psd_fpga_top.vh"
    
// ***********************************************************
// Include local parameters definitions for the GPIO ports
// DO NOT modify!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!
// It is auto-generated by the assign_gpio.tcl generator
// ***********************************************************

`include    "gpio_defines.vh"

// Define a bunch of wires
// Hand generated but include reduces clutter in this file

`include    "psd_fpga_top_wires.vh"

// $$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$

// *********************************     
// Instaniate the ublaze wrapper
// *********************************    
 
    psd_ublaze_wrapper  u0(
        .clk10(clk10),
        .gpio0_in(gpio0_in),
        .gpio0_out(gpio0_out),
        .gpio1_in(gpio1_in),
        .gpio1_out(gpio1_out),
        .gpio2_in(gpio2_in),
        .gpio2_out(gpio2_out),
        .gpio3_in(gpio3_in),
        .gpio3_out(gpio3_out),
        .iic_rtl_0_scl_io(i2c_scl),
        .iic_rtl_0_sda_io(i2c_sda),
        .mclk(mclk),
        .reset(ublaze_reset),
        .sys_clk(sys_clk),
        .uart_rtl_1_baudoutn(baudout),
        .uart_rtl_1_ctsn(cts),
        .uart_rtl_1_dcdn(dcd),
        .uart_rtl_1_ddis(ddis),
        .uart_rtl_1_dsrn(dsr),
        .uart_rtl_1_dtrn(dtr),
        .uart_rtl_1_out1n(out1),
        .uart_rtl_1_out2n(out2),
        .uart_rtl_1_ri(ri),
        .uart_rtl_1_rtsn(rts),
        .uart_rtl_1_rxd(uart_rx),
        .uart_rtl_1_rxrdyn(rxrdy),
        .uart_rtl_1_txd(uart_tx),
        .uart_rtl_1_txrdyn(txrdy),
        .fifo_data(fifo_data),
        .tlast(tlast),
        .tready(tready),
        .tvalid(tvalid)
    ) ;

// ********************************************************  
// Instantiate the custom block
// mclk is 100 MHz clock from ublaze
//
// GPIO ports 2 and 3 are for the exclusive use of uBlaze
// **********************************************************

    psd_custom_block u1(
        .mclk(mclk) ,
        .mrst(custom_block_reset) ,
        .led(led) ,
        .gpio0_in(gpio0_in) ,
        .gpio1_in(gpio1_in) ,
        .gpio0_out(gpio0_out) ,
        .gpio1_out(gpio1_out) ,         
        .tready(tready) ,
        .adc_sdo(adc_sdo) ,
        .adc_sclk(adc_sclk) ,
        .adc_conv(adc_conv) ,
        .fifo_data(fifo_data) ,
        .tlast(tlast) ,
        .tvalid(tvalid) ,
        .common_stop(common_stop)        
    ) ;

// ********************************    
// Assign of pins to signals
// **********************************

// Reset stuff

    assign  ublaze_reset = dummy_reset ;
    assign  custom_block_reset = dummy_reset ;

// Make some connections for the UART

    assign dcd = 1'b1 ;
    assign dsr = 1'b1 ;
//    assign dsr = dtr ;
    assign ri = 1'b1 ;
    assign cts = rts ;
    
// Make connections for the ADCs 
   
    assign  adc_sclk_0 = adc_sclk[0] ;
    assign  conv_0 = adc_conv[0] ;

    assign  adc_sdo[0] = 1'b0 ;     // PSD 0 Sub-Channel A
    assign  adc_sdo[1] = 1'b0 ;     // PSD 0 Sub-Channel B    
    assign  adc_sdo[2] = 1'b0 ;     // PSD 0 Sub-Channel C   
    assign  adc_sdo[3] = sdo_t_0 ;  // PSD 0 Sub-Channel T
    assign  adc_sdo[4] = 1'b0 ;     // PSD 1 Sub-Channel A    
    assign  adc_sdo[5] = 1'b0 ;     // PSD 1 Sub-Channel B     
    assign  adc_sdo[6] = 1'b0 ;     // PSD 1 Sub-Channel C  
    assign  adc_sdo[7] = 1'b0 ;     // PSD 1 Sub-Channel T 
    
// Timestamp related stuff
// This is just a place keeper

    assign  tstamp_clk = clk10 ;
    assign  tstamp_rst = 1'b0 ;
    
// *****************************************************
// The gpio_assigns.h file AUTO-GENERATED
// NEVER DIRECTLY MODIFY IT!!!!
// *****************************************************

`include "gpio_assigns.vh"

// *****************************************************
// Create bi-directional cfd_ad bus
// *****************************************************
   
    assign  cfd_ad[7:0] = cfd_write ? cfd_ad_out[7:0] : 8'bzzzz_zzzz ;
    assign  cfd_ad_in[7:0] = cfd_ad[7:0] ;
    
// *****************************************************
// TEMP:   Create PSD0 test intx output to be routed out to backboard.
// TODO: Implement a mux for this in custom block. 
// *****************************************************  
    
 assign intx_out =  psd_intx_out_0; 
    
    
// assign or_connect = cfd_or_connect;
//assign cfd_or_connect = cfd_or ;

endmodule
