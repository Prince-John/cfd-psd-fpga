`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07/25/2024 04:32:57 PM
// Design Name: 
// Module Name: psd_custom_block
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
// In this version of the custom block, we will test out the AXI Stream FIFO
// by streaming ADC7687 adc data to it!
// So we are also testing out the ADC register and associated control
//
// FIFO data is 32 bits wide :
//      Upper byte is a tag or data type indentifier
//      Lower 3 bytes are to be used for data
//
// The gpios are ALL inputs to the custom block here
//
//////////////////////////////////////////////////////////////////////////////////

module psd_custom_block(

    input   mclk ,
    input   mrst ,
    output  [1:0] led ,
    input   [31:0] gpio0_in ,
    input   [31:0] gpio1_in ,   
    output  [31:0] gpio0_out ,
    output  [31:0] gpio1_out ,      
    input   tready ,
    input   [7:0] adc_sdo ,
    output  [1:0] adc_sclk ,
    output  [1:0] adc_conv ,
    output  [31:0] fifo_data ,
    output  tlast ,
    output  tvalid ,
    input   common_stop 
    
   ) ;
   
// ***********************************************************
// Include local parameters definitions for the GPIO ports
// DO NOT modify!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!
// It is auto-generated by the assign_gpio.tcl generator
// ***********************************************************

`include    "gpio_defines.vh"

    
// ***************************    
// Wire up the input ports
// ***************************

    wire    [7:0] p0_in ;
    wire    [7:0] p1_in ;    
    wire    [7:0] p2_in ;    
    wire    [7:0] p3_in ;  
    wire    [7:0] p4_in ;
    wire    [7:0] p5_in ;    
    wire    [7:0] p6_in ;    
    wire    [7:0] p7_in ; 

    assign  p0_in[0] = tready ;
    assign  p0_in[7:1] = 7'd0 ;
    
    assign  p1_in[5:0] = gpio0_in[BOARD_ID_5 : BOARD_ID_0] ;
    assign  p1_in[7:6] = 2'd0 ;
    
    assign  p2_in[7:0] = 8'd0 ;        
    assign  p3_in[7:0] = 8'd0 ;  
    assign  p4_in[7:0] = 8'd0 ;     
    assign  p5_in[7:0] = 8'd0 ;     
    assign  p6_in[7:0] = 8'd0 ;     
    assign  p7_in[7:0] = 8'd0 ;     
       
    
// *******************************
// Wire up the output ports
// *******************************
      
    wire    [7:0] p0_out ;
    wire    [7:0] p1_out ;    
    wire    [7:0] p2_out ;
    wire    [7:0] p3_out ;
    wire    [7:0] p4_out ;
    wire    [7:0] p5_out ;    
    wire    [7:0] p6_out ;
    wire    [7:0] p7_out ;  
     
// ^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^  
//  OUTPUT PORT 0
// Picoblaze will use it as a heartbeat indicator
// ^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^

    assign  led[0] = p0_out[0] ;
    assign  led[1] = p0_out[1] ;
    
// ^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^  
//  OUTPUT PORT 1
//  Assign adc clocks and conv signals to port bits!!!
// ^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^
 
    assign  adc_sclk[0] = p1_out[0] ;
    assign  adc_sclk[1] = p1_out[1] ;
    assign  adc_conv[0] = p1_out[2] ; 
    assign  adc_conv[1] = p1_out[3] ;
 
// Use 3 bits to select which ADC should drive the fifo data bus
   
    wire    [2:0] adc_mux_sel ;
    wire    adc_reg_reset ;
    
    assign  adc_mux_sel = p1_out[6:4] ; 
    assign  adc_reg_reset = p1_out[7] ;

// ^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^  
//  OUTPUT PORT 2
// Use output port 2 to put out data type identifier
// ^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^
   
    wire    [7:0] data_id ;
    assign  data_id = p2_out ;
    
// ^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^  
//  OUTPUT PORT 3
//  Byte going out to tdc_reg
// ^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^    
    
    wire    [7:0] tdc_byte ;
    assign  tdc_byte = p3_out ;
    
// ^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^  
//  OUTPUT PORT 4
//  Byte going out to tdc_reg
// ^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^ 
    
    wire    [2:0] tdc_reg_ld ;
    assign  tdc_reg_ld = p4_out[2:0] ;
    
    wire    tdc_reg_rst, tdc_reg_shift ;
    assign  tdc_reg_rst = p4_out[3] ;
    assign  tdc_reg_shift = p4_out[4] ;
    assign  tdc_sclk = p4_out[5] ;
    
// $$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$
// Instantiate our Picoblaze 6 microcontroller
// $$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$  
     
    picoblaze_controller  proc0 (
            .clk(mclk),
            .reset(mrst),
            .P0_in(p0_in),
            .P1_in(p1_in),
            .P2_in(p2_in),
            .P3_in(p3_in),  
            .P4_in(p4_in),
            .P5_in(p5_in),
            .P6_in(p6_in),
            .P7_in(p7_in),                             
            .P0_out(p0_out),
            .P1_out(p1_out),
            .P2_out(p2_out),
            .P3_out(p3_out),
            .P4_out(p4_out),
            .P5_out(p5_out),
            .P6_out(p6_out),
            .P7_out(p7_out),                        
            .tvalid(tvalid),
            .tlast(tlast)        
    ) ;
    
// **************************************************************
// Insert a bank of 4 ADC registers for PSD chip 0
// They perform serial-to-parallel conversion
// Asynchronous reset that picoblaze can use to clear register
// ************************************************************

    reg     [15:0] adc_0_reg_a ;
    reg     [15:0] adc_0_reg_b ;    
    reg     [15:0] adc_0_reg_c ;
    reg     [15:0] adc_0_reg_t ;    
    
    always @(negedge adc_sclk[0] or posedge adc_reg_reset) begin
        if (adc_reg_reset) begin
            adc_0_reg_a <= 16'd0 ;
            adc_0_reg_b <= 16'd0 ;
            adc_0_reg_c <= 16'd0 ;
            adc_0_reg_t <= 16'd0 ;            
        end else begin
            adc_0_reg_a <= {adc_0_reg_a[14:0], adc_sdo[0]} ;
            adc_0_reg_b <= {adc_0_reg_b[14:0], adc_sdo[1]} ;           
            adc_0_reg_c <= {adc_0_reg_c[14:0], adc_sdo[2]} ;            
            adc_0_reg_t <= {adc_0_reg_t[14:0], adc_sdo[3]} ;            
        end        
	end
    
// *********************************************************
// Insert a bank of 4 ADC registers for PSD chip 1
// They perform serial-to-parallel conversion
// *********************************************************

    reg     [15:0] adc_1_reg_a ;
    reg     [15:0] adc_1_reg_b ;    
    reg     [15:0] adc_1_reg_c ;
    reg     [15:0] adc_1_reg_t ;    
    
    always @(negedge adc_sclk[1] or posedge adc_reg_reset) begin
        if (adc_reg_reset) begin
            adc_1_reg_a <= 16'd0 ;
            adc_1_reg_b <= 16'd0 ;
            adc_1_reg_c <= 16'd0 ;
            adc_1_reg_t <= 16'd0 ;            
        end else begin
            adc_1_reg_a <= {adc_1_reg_a[14:0], adc_sdo[4]} ;
            adc_1_reg_b <= {adc_1_reg_b[14:0], adc_sdo[5]} ;           
            adc_1_reg_c <= {adc_1_reg_c[14:0], adc_sdo[6]} ;            
            adc_1_reg_t <= {adc_1_reg_t[14:0], adc_sdo[7]} ;            
        end        
	end   
	
// **************************************************************
// Implement a MUX to pick what drives the fifo data bus
// Bits 2-4 will select which ADC reg drive fifo
// Port 2 will be the data tag identifier
// **************************************************************

    reg    [31:0] adc_reg ;
    always @(*) begin   
        case (adc_mux_sel)
            3'd0:   adc_reg = {data_id, 8'd0, adc_0_reg_a} ;
            3'd1:   adc_reg = {data_id, 8'd0, adc_0_reg_b} ;       
            3'd2:   adc_reg = {data_id, 8'd0, adc_0_reg_c} ;        
            3'd3:   adc_reg = {data_id, 8'd0, adc_0_reg_t} ;
            3'd4:   adc_reg = {data_id, 8'd0, adc_1_reg_a} ;
            3'd5:   adc_reg = {data_id, 8'd0, adc_1_reg_b} ;       
            3'd6:   adc_reg = {data_id, 8'd0, adc_1_reg_c} ;        
            3'd7:   adc_reg = {data_id, 8'd0, adc_1_reg_t} ;
        endcase
    end   
    

// ************************************************

    assign  fifo_data = adc_reg ;
    
endmodule