../gpio/gpio_defines.vh